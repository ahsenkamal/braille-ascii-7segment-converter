module BrailleTo7Segment(i,o1,o0);

input [1:6]i;
output [1:7]o1,o0;

assign o1[1] = (i[1]&(~i[6])) | (i[4]&(~i[5])) | (i[1]&i[2]) | ((~i[2])&i[5]&(~i[6])) | (i[3]&(~i[4])&i[6]) | (i[1]&(~i[3])&i[5]) | (i[2]&i[3]&(~i[6])) | ((~i[3])&(~i[5])&(~i[6])) | (i[2]&(~i[3])&i[4]) | ((~i[1])&(~i[2])&i[3]&i[6]); 
assign o1[2] = ((~i[3])&(~i[4])&i[6]) | (i[2]&i[3]&(~i[6])) | ((~i[3])&i[5]&i[6]) | (i[2]&i[3]&(~i[5])) | (i[2]&(~i[4])&i[5]) | ((~i[1])&i[2]&i[6]) | (i[1]&(~i[2])&i[3]&i[5]) | (i[1]&(~i[2])&i[3]&i[4]) | (i[1]&i[2]&i[4]&(~i[6])) | (i[3]&(~i[4])&(~i[5])&(~i[6])) | ((~i[1])&(~i[2])&(~i[3])&(~i[4])) | ((~i[1])&(~i[3])&i[4]&(~i[5])&(~i[6]));
assign o1[3] = 1;
assign o1[4] = (i[4]&(~i[5])&i[6]) | ((~i[2])&(~i[3])&(~i[6])) | (i[1]&i[2]&i[6]) | (i[3]&(~i[4])&i[6]) | ((~i[3])&(~i[4])&(~i[5])&(~i[6])) | (i[1]&(~i[3])&i[5]&i[6]) | ((~i[1])&i[2]&(~i[3])&i[4]) | ((~i[1])&i[3]&i[5]&(~i[6])) | (i[1]&i[2]&i[3]&i[4]) | ((~i[1])&(~i[2])&i[3]&i[4]) | (i[1]&i[2]&i[3]&i[5]);
assign o1[5] = (i[2]&i[3]&i[5]&(~i[6])) | (i[1]&(~i[2])&(~i[3])&(~i[6])) | (i[2]&(~i[3])&(~i[4])&(~i[5])&(~i[6])) | ((~i[1])&i[2]&i[4]&i[5]&(~i[6])) | (i[1]&(~i[3])&(~i[4])&i[5]&i[6]) | (i[1]&i[3]&(~i[4])&(~i[5])&i[6]) | (i[1]&i[2]&(~i[3])&i[4]&i[6]) | (i[1]&i[2]&i[4]&i[5]&i[6]) | (i[1]&i[2]&i[3]&i[4]&(~i[6])) | ((~i[1])&i[2]&i[3]&i[4]&(~i[5])&i[6]);
assign o1[6] = ((~i[2])&i[6]) | (i[3]&i[4]&i[6]) | (i[3]&(~i[5])&i[6]) | ((~i[1])&(~i[2])&i[3]) | ((~i[1])&(~i[5])&i[6]) | (i[1]&i[4]&i[6]) | (i[1]&(~i[2])&(~i[3])) | ((~i[1])&i[4]&i[5]&(~i[6])) | (i[1]&i[2]&i[3]&i[4]) | ((~i[3])&(~i[4])&i[5]&i[6]) | ((~i[1])&i[2]&(~i[3])&(~i[6])) | (i[2]&i[3]&i[5]&(~i[6])) | (i[1]&(~i[3])&(~i[4])&(~i[5])&(~i[6]));
assign o1[7] = (i[6]) | ((~i[1])&(~i[2])) | ((~i[1])&(~i[3])) | ((~i[2])&(~i[3])) | ((~i[3])&(~i[4])&(~i[5])) | (i[2]&i[3]&i[5]) | (i[1]&i[2]&i[3]&i[4]);

assign o0[1] = (i[1]&(~i[2])) | ((~i[4])&i[5]) | (i[1]&(~i[5])) | (i[2]&(~i[3])&i[6]) | ((~i[2])&i[3]&i[6]) | ((~i[2])&(~i[4])&(~i[6])) | (i[4]&(~i[5])&i[6]) | ((~i[1])&(~i[3])&i[5]) | (i[3]&(~i[4])&(~i[6]));
assign o0[2] = ((~i[1])&(~i[6])) | (i[5]&(~i[6])) | (i[1]&i[4]) | ((~i[2])&(~i[5])&i[6]) | ((~i[2])&(~i[3])&i[4]) | (i[2]&(~i[4])&i[5]) | ((~i[1])&i[2]&i[3]) | (i[1]&i[3]&i[5]) | (i[1]&(~i[3])&(~i[5])&i[6]);
assign o0[3] = (i[5]&i[6]) | (i[2]&(~i[5])) | ((~i[1])&(~i[3])&i[6]) | ((~i[1])&(~i[4])&i[5]) | ((~i[2])&(~i[3])&i[4]) | ((~i[2])&i[3]&(~i[4])) | (i[3]&i[4]&(~i[6])) | (i[1]&(~i[2])&(~i[6])) | (i[1]&(~i[3])&i[4]);
assign o0[4] = ((~i[4])&i[5]&i[6]) | ((~i[3])&i[4]&i[6]) | (i[1]&(~i[2])&(~i[4])) | (i[3]&(~i[4])&(~i[6])) | (i[1]&i[3]&(~i[4])) | ((~i[2])&i[3]&i[6]) | ((~i[2])&(~i[4])&(~i[6])) | (i[1]&(~i[4])&(~i[6])) | (i[1]&(~i[2])&i[5]) | (i[1]&i[2]&i[4]&(~i[5])) | ((~i[1])&i[2]&(~i[3])&i[6]) | ((~i[1])&i[2]&(~i[3])&i[4]&i[5]);
assign o0[5] = (i[1]&(~i[2])&(~i[5])&i[6]) | (i[1]&(~i[2])&i[4]&i[5]) | (i[1]&i[3]&(~i[4])&i[6]) | (i[1]&i[2]&(~i[5])&(~i[6])) | (i[1]&i[2]&(~i[4])&i[5]) | ((~i[2])&(~i[3])&i[4]&i[5]&i[6]) | ((~i[1])&(~i[2])&i[3]&(~i[4])&i[5]) | ((~i[2])&i[3]&i[4]&(~i[5])&i[6]) | ((~i[1])&(~i[2])&(~i[3])&(~i[4])&(~i[5])&(~i[6])) | ((~i[1])&i[2]&(~i[3])&(~i[4])&(~i[5])&i[6]) | ((~i[1])&i[2]&(~i[3])&i[4]&i[5]&(~i[6]));
assign o0[6] = ((~i[2])&(~i[4])&i[5]) | ((~i[2])&i[5]&i[6]) | (i[1]&(~i[2])&i[5]) | ((~i[1])&(~i[3])&(~i[5])&i[6]) | ((~i[1])&(~i[3])&i[4]&(~i[5])) | ((~i[2])&(~i[3])&i[4]&i[6]) | ((~i[3])&i[4]&i[5]&i[6]) | ((~i[2])&i[3]&(~i[4])&(~i[6])) | (i[2]&(~i[3])&(~i[5])&(~i[6])) | (i[2]&i[4]&(~i[5])&(~i[6])) | (i[1]&(~i[2])&(~i[4])&(~i[6])) | (i[1]&(~i[4])&i[5]&i[6]) | (i[1]&i[3]&(~i[4])&(~i[5])) | ((~i[1])&i[3]&i[4]&i[5]&(~i[6]));
assign o0[7] = ((~i[1])&(~i[2])&i[6]) | ((~i[4])&(~i[5])&(~i[6])) | ((~i[1])&(~i[3])&(~i[5])) | (i[1]&(~i[4])&(~i[6])) | ((~i[2])&(~i[3])&(~i[4])) | (i[1]&(~i[2])&i[5]&(~i[6])) | (i[2]&i[3]&(~i[4])&i[5]) | (i[1]&i[4]&(~i[5])&i[6]) | ((~i[1])&i[2]&i[4]&(~i[6])) | (i[2]&(~i[3])&i[5]&i[6]) | (i[1]&i[2]&i[3]&(~i[4])) | ((~i[2])&i[3]&i[4]&i[5]&(~i[6]));

endmodule